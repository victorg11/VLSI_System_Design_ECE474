class input_data;
rand bit[31:0] dataA;
rand bit[31:0] dataB;

// constraint positive {dataA > 0}; //values must be positive
// constraint positive {dataB >= 0}; //values must be positive

endclass
